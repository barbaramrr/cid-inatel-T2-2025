module not_gate (
    output b,
    input a
);

    not (b,a);

endmodule